module RAM_512x16_clarinet (
    input [8:0] ram_addr,
    input [15:0] ram_wdata,
    output [15:0] ram_rdata,
    input ce,
    input clk,
    input we,
    input re);

    wire [15:0] ram_rdata0;
    wire [15:0] ram_rdata1;

    assign ram_rdata = ram_addr[8] ? ram_rdata1 : ram_rdata0;

    SB_RAM40_4K RAM_inst0(
        .RDATA(ram_rdata0),
        .RADDR({3'b000,ram_addr[7:0]}),
        .RCLK(clk),
        .RCLKE(re&ce),
        .RE(re&ce),
        .WDATA(ram_wdata),
        .WADDR({3'b000,ram_addr[7:0]}),
        .WCLK(clk),
        .WCLKE(we&ce),
        .WE(we&ce),
        .MASK(16'h0000));
    defparam RAM_inst0.READ_MODE =0;
    defparam RAM_inst0.WRITE_MODE =0;

    SB_RAM40_4K RAM_inst1(
        .RDATA(ram_rdata1),
        .RADDR({3'b000,ram_addr[7:0]}),
        .RCLK(clk),
        .RCLKE(re&ce),
        .RE(re&ce),
        .WDATA(ram_wdata),
        .WADDR({3'b000,ram_addr[7:0]}),
        .WCLK(clk),
        .WCLKE(we&ce),
        .WE(we&ce),
        .MASK(16'h0000));
    defparam RAM_inst0.READ_MODE =0;
    defparam RAM_inst0.WRITE_MODE =0;

    /*clarinet */
    defparam RAM_inst0.INIT_0 = 256'h7C19_75E6_6F9F_695A_6332_5D3C_578C_5231_4D39_48AB_448C_40DE_3D9C_3AC1_3845_361E;
    defparam RAM_inst0.INIT_1 = 256'hA734_A777_A78C_A764_A6ED_A618_A4D5_A317_A0D2_9E01_9A9F_96AF_9237_8D41_87DE_821E;
    defparam RAM_inst0.INIT_2 = 256'h97CA_9989_9B3A_9CD0_9E43_9F8F_A0B2_A1B0_A28E_A352_A402_A4A5_A53E_A5CF_A657_A6D0;
    defparam RAM_inst0.INIT_3 = 256'hAD2A_A88B_A3FF_9FB1_9BC5_985A_9585_9356_91D1_90F4_90B6_9105_91CD_92F8_946B_960E;
    defparam RAM_inst0.INIT_4 = 256'h9B7F_A1EE_A82D_AE0C_B35D_B7F6_BBB3_BE79_C035_C0E0_C07C_BF17_BCC6_B9A9_B5E8_B1AE;
    defparam RAM_inst0.INIT_5 = 256'h721E_7120_704D_6FBE_6F8A_6FC8_7090_71F5_7406_76CE_7A4F_7E86_8367_88DC_8ECA_950E;
    defparam RAM_inst0.INIT_6 = 256'h7CE4_7C51_7BD6_7B6B_7B0A_7AAD_7A4D_79E2_7965_78D1_7822_7755_766B_7568_7453_7335;
    defparam RAM_inst0.INIT_7 = 256'h9058_8F86_8E79_8D3B_8BD7_8A59_88CD_873C_85B2_8436_82CF_8182_8055_7F48_7E5C_7D91;
    defparam RAM_inst0.INIT_8 = 256'h8889_87EF_87CB_8813_88B5_899E_8ABA_8BF1_8D2D_8E5A_8F64_903B_90D4_9126_912C_90E7;
    defparam RAM_inst0.INIT_9 = 256'hB4DF_B30B_B0CD_AE2B_AB30_A7EA_A46C_A0CA_9D1C_997B_95FF_92C1_8FD5_8D4E_8B3A_89A1;
    defparam RAM_inst0.INIT_A = 256'hA579_A80F_AA82_ACCE_AEEF_B0E1_B2A2_B42D_B57E_B68F_B75C_B7DB_B807_B7D6_B743_B647;
    defparam RAM_inst0.INIT_B = 256'h8D50_8C0A_8B40_8AF4_8B27_8BD4_8CF4_8E7D_9062_9294_9505_97A5_9A63_9D31_A001_A2C7;
    defparam RAM_inst0.INIT_C = 256'hC671_C246_BE11_B9D6_B59B_B164_AD36_A91A_A515_A133_9D7C_99FC_96BE_93D0_913C_8F0E;
    defparam RAM_inst0.INIT_D = 256'hF776_F5AA_F3B6_F199_EF50_ECD7_EA2F_E755_E44A_E110_DDA9_DA18_D662_D28B_CE98_CA8E;
    defparam RAM_inst0.INIT_E = 256'hF258_F5F6_F8FF_FB73_FD56_FEB0_FF8C_FFF7_FFFE_FFB0_FF17_FE42_FD37_FC00_FAA2_F91E;
    defparam RAM_inst0.INIT_F = 256'h975D_9C3E_A164_A6D1_AC86_B27D_B8AD_BF08_C57D_CBF6_D25D_D899_DE94_E437_E96D_EE27;

    defparam RAM_inst1.INIT_0 = 256'h55C7_5904_5C99_6070_6477_689D_6CD1_7109_753C_7966_7D89_81A8_85CA_89FB_8E47_92B9;
    defparam RAM_inst1.INIT_1 = 256'h62E8_6001_5D08_5A11_5732_5484_521C_5012_4E77_4D5F_4CD4_4CE0_4D86_4EC6_5098_52F2;
    defparam RAM_inst1.INIT_2 = 256'h7602_758D_7525_74C6_7466_73FD_737F_72E2_721A_711D_6FE3_6E64_6C9E_6A90_683D_65AC;
    defparam RAM_inst1.INIT_3 = 256'h7E47_7E8C_7EA1_7E87_7E40_7DD3_7D43_7C97_7BD6_7B07_7A33_795F_7892_77D3_7724_7689;
    defparam RAM_inst1.INIT_4 = 256'h699E_6ADF_6C44_6DC5_6F5B_70FD_72A4_7448_75E1_7768_78D6_7A25_7B50_7C53_7D29_7DD1;
    defparam RAM_inst1.INIT_5 = 256'h6E5D_6D52_6C3E_6B27_6A18_6919_6833_676F_66D5_666B_6636_663A_6678_66F1_67A2_6888;
    defparam RAM_inst1.INIT_6 = 256'h763D_75C4_7558_74FB_74A9_745F_741B_73D6_738A_7334_72CC_724F_71B9_7108_703C_6F58;
    defparam RAM_inst1.INIT_7 = 256'h8027_7F81_7EDC_7E3B_7D9D_7D01_7C65_7BC8_7B29_7A86_79E1_793B_7895_77F3_7757_76C4;
    defparam RAM_inst1.INIT_8 = 256'h6FE7_73B0_771E_7A22_7CB3_7ECC_806E_819E_8266_82D1_82EE_82CA_8275_81FC_816B_80CC;
    defparam RAM_inst1.INIT_9 = 256'h511F_4F02_4D61_4C52_4BE4_4C24_4D14_4EB4_50F9_53D6_5735_5AFC_5F10_634F_679D_6BD9;
    defparam RAM_inst1.INIT_A = 256'h72CC_723F_7181_708B_6F58_6DE2_6C24_6A1E_67D0_6540_6278_5F84_5C78_5968_566D_53A1;
    defparam RAM_inst1.INIT_B = 256'h61E6_64BC_6755_69AD_6BC0_6D8C_6F14_7059_715F_722A_72C1_7328_7364_7378_7366_732D;
    defparam RAM_inst1.INIT_C = 256'h2C35_2EF6_31E7_3502_3841_3B9E_3F15_42A1_463B_49DF_4D85_5126_54BB_583B_5B9D_5ED9;
    defparam RAM_inst1.INIT_D = 256'h2766_25DE_2465_230C_21E2_20F5_2050_1FFC_1FFF_205D_2118_222C_2398_2555_275E_29AB;
    defparam RAM_inst1.INIT_E = 256'h2C0B_2C98_2D31_2DCC_2E5D_2ED9_2F33_2F62_2F5C_2F1C_2E9E_2DE1_2CE9_2BBC_2A64_28EE;
    defparam RAM_inst1.INIT_F = 256'h3442_32A6_3141_3009_2EF8_2E0A_2D39_2C86_2BF1_2B7A_2B25_2AF2_2AE4_2AFB_2B36_2B92;

endmodule
