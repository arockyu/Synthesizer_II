/************************************************************************
* Extended Hex to 7-Seg decoder unit
*
*************************************************************************
* input  oe            : LED patter outoput enable (Active-High)
* input [4:0] hex      : 1 digit hex(4-bit) input
* output [6:0] pat7seg : coded 7seg pattern output {g,f,e,d,c,b,a}
***************************************************************************
*  
* 
****************************************************************************/

module hexto7seg_ex(
    input oe,
    input [4:0] hex,
    output [6:0] pat7seg);

    assign pat7seg = ( oe  ==  1'b0  ) ? 7'b0000000 : 
                     ( hex ==  5'h00 ) ? 7'b0111111 :
                     ( hex ==  5'h01 ) ? 7'b0000110 :     
                     ( hex ==  5'h02 ) ? 7'b1011011 :     
                     ( hex ==  5'h03 ) ? 7'b1001111 : 
                     ( hex ==  5'h04 ) ? 7'b1100110 : 
                     ( hex ==  5'h05 ) ? 7'b1101101 : 
                     ( hex ==  5'h06 ) ? 7'b1111101 : 
                     ( hex ==  5'h07 ) ? 7'b0000111 : 
                     ( hex ==  5'h08 ) ? 7'b1111111 : 
                     ( hex ==  5'h09 ) ? 7'b1101111 : 
                     ( hex ==  5'h0a ) ? 7'b1110111 : //a
                     ( hex ==  5'h0b ) ? 7'b1111100 : //b
                     ( hex ==  5'h0c ) ? 7'b0111001 : //c
                     ( hex ==  5'h0d ) ? 7'b1011110 : //d
                     ( hex ==  5'h0e ) ? 7'b1111001 : //e
                     ( hex ==  5'h0f ) ? 7'b1110001 : //f
                     ( hex ==  5'h10 ) ? 7'b0111101 : //G
                     ( hex ==  5'h11 ) ? 7'b1000000 : //-
                     ( hex ==  5'h12 ) ? 7'b1011100 : //o                   
                     ( hex ==  5'h13 ) ? 7'b0111000 : //L
                     ( hex ==  5'h14 ) ? 7'b1010000 : //r
                     ( hex ==  5'h15 ) ? 7'b1010100 : 7'b0000000;  //n                
endmodule