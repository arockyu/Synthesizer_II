module RAM_512x16_trum (
    input [8:0] ram_addr,
    input [15:0] ram_wdata,
    output [15:0] ram_rdata,
    input ce,
    input clk,
    input we,
    input re);

    wire [15:0] ram_rdata0;
    wire [15:0] ram_rdata1;

    assign ram_rdata = ram_addr[8] ? ram_rdata1 : ram_rdata0;

    SB_RAM40_4K RAM_inst0(
        .RDATA(ram_rdata0),
        .RADDR({3'b000,ram_addr[7:0]}),
        .RCLK(clk),
        .RCLKE(re&ce),
        .RE(re&ce),
        .WDATA(ram_wdata),
        .WADDR({3'b000,ram_addr[7:0]}),
        .WCLK(clk),
        .WCLKE(we&ce),
        .WE(we&ce),
        .MASK(16'h0000));
    defparam RAM_inst0.READ_MODE =0;
    defparam RAM_inst0.WRITE_MODE =0;

    SB_RAM40_4K RAM_inst1(
        .RDATA(ram_rdata1),
        .RADDR({3'b000,ram_addr[7:0]}),
        .RCLK(clk),
        .RCLKE(re&ce),
        .RE(re&ce),
        .WDATA(ram_wdata),
        .WADDR({3'b000,ram_addr[7:0]}),
        .WCLK(clk),
        .WCLKE(we&ce),
        .WE(we&ce),
        .MASK(16'h0000));
    defparam RAM_inst0.READ_MODE =0;
    defparam RAM_inst0.WRITE_MODE =0;

    /*trumpet*/
    defparam RAM_inst0.INIT_0 = 256'h882C_8606_841F_8276_8104_7FBD_7E94_7D7C_7C68_7B55_7A3F_792A_7820_772B_7658_75B0;
    defparam RAM_inst0.INIT_1 = 256'hB13F_ABFB_A7CD_A492_A213_A018_9E65_9CC8_9B17_9937_971D_94C9_9248_8FAD_8D10_8A89;
    defparam RAM_inst0.INIT_2 = 256'hDCA4_E8D2_F2BD_FA07_FE77_FFFE_FEB6_FADF_F4D9_ED1F_E438_DAB1_D10F_C7C9_BF3D_B7AD;
    defparam RAM_inst0.INIT_3 = 256'h4BF0_4BE0_4C7D_4DFF_50A3_54A7_5A42_619F_6AD4_75DE_8299_90C2_9FF7_AFBE_BF84_CEAF;
    defparam RAM_inst0.INIT_4 = 256'h7166_6F53_6CBA_69B9_6672_630C_5FA9_5C68_5962_56A4_5437_5218_5046_4EBB_4D77_4C82;
    defparam RAM_inst0.INIT_5 = 256'h6D00_6C3F_6BB3_6B6E_6B7C_6BE4_6CA4_6DAF_6EF2_704F_71A3_72C7_7396_73EE_73B7_72E0;
    defparam RAM_inst0.INIT_6 = 256'h7C57_7B4F_7A35_7916_77FC_76F0_75F5_750C_7430_735C_7287_71AC_70C5_6FD3_6EDA_6DE5;
    defparam RAM_inst0.INIT_7 = 256'h7F25_7EBE_7E67_7E2B_7E0F_7E13_7E34_7E6A_7EA9_7EE3_7F09_7F0E_7EE7_7E8D_7DFF_7D3F;
    defparam RAM_inst0.INIT_8 = 256'h80C5_805B_800A_7FD8_7FC6_7FD2_7FF7_8029_805F_808C_80A7_80A7_8089_804D_7FF8_7F92;
    defparam RAM_inst0.INIT_9 = 256'h801C_8063_80B6_8115_817D_81E8_824D_82A5_82E5_8307_8305_82E0_8298_8234_81BD_813F;
    defparam RAM_inst0.INIT_A = 256'h79F3_7A0A_7A46_7AA3_7B1D_7BAB_7C45_7CE2_7D78_7E00_7E77_7ED9_7F2A_7F6C_7FA6_7FDF;
    defparam RAM_inst0.INIT_B = 256'h7D07_7CE6_7CCD_7CBA_7CA7_7C92_7C74_7C4A_7C11_7BCA_7B76_7B1B_7AC0_7A6C_7A29_79FE;
    defparam RAM_inst0.INIT_C = 256'h7B79_7BBE_7C13_7C71_7CD2_7D2F_7D7F_7DBE_7DE7_7DFA_7DF6_7DE0_7DBB_7D8D_7D5D_7D2F;
    defparam RAM_inst0.INIT_D = 256'h7F48_7EB7_7E35_7DC2_7D5D_7D01_7CAC_7C5D_7C13_7BCE_7B91_7B5F_7B3B_7B2A_7B2E_7B48;
    defparam RAM_inst0.INIT_E = 256'h80A5_8177_823B_82E7_8374_83D8_8411_841A_83F4_83A3_832E_829B_81F5_8145_8093_7FE8;
    defparam RAM_inst0.INIT_F = 256'h7996_7981_7987_79A5_79D7_7A1A_7A6B_7AC9_7B34_7BAD_7C35_7CCE_7D78_7E33_7EFC_7FCF;

    defparam RAM_inst1.INIT_0 = 256'h7F93_7FB7_7FC8_7FBE_7F95_7F4C_7EE2_7E5B_7DBD_7D12_7C61_7BB4_7B15_7A8B_7A1B_79C9;
    defparam RAM_inst1.INIT_1 = 256'h81C4_815C_80FA_809A_803E_7FE6_7F95_7F4D_7F13_7EE9_7ED3_7ED1_7EE2_7F04_7F32_7F64;
    defparam RAM_inst1.INIT_2 = 256'h8813_883E_884A_8835_87FE_87A7_8736_86B0_861A_857D_84DE_8443_83AF_8326_82A6_8231;
    defparam RAM_inst1.INIT_3 = 256'h7FEB_8087_8120_81B4_8242_82CD_8353_83D9_845F_84E6_856E_85F6_867B_86F9_876B_87CA;
    defparam RAM_inst1.INIT_4 = 256'h7B9E_7BA8_7BAF_7BB7_7BBF_7BCC_7BE0_7C00_7C2F_7C6F_7CC2_7D27_7D9F_7E25_7EB6_7F4F;
    defparam RAM_inst1.INIT_5 = 256'h7B36_7B64_7B87_7B9F_7BAA_7BAB_7BA4_7B98_7B8B_7B7F_7B77_7B75_7B77_7B7E_7B88_7B93;
    defparam RAM_inst1.INIT_6 = 256'h7CC6_7C89_7C3E_7BE9_7B8E_7B33_7AE0_7A9A_7A65_7A45_7A3C_7A48_7A66_7A93_7AC8_7B00;
    defparam RAM_inst1.INIT_7 = 256'h7CB3_7CDC_7CF7_7D05_7D0B_7D0B_7D08_7D07_7D09_7D0E_7D15_7D1D_7D21_7D1E_7D0F_7CF3;
    defparam RAM_inst1.INIT_8 = 256'h7C51_7C08_7BBB_7B71_7B2E_7AF7_7AD3_7AC4_7ACB_7AE9_7B1A_7B5B_7BA4_7BF1_7C3B_7C7D;
    defparam RAM_inst1.INIT_9 = 256'h8162_8108_809B_8022_7FA6_7F2D_7EBD_7E5A_7E07_7DC3_7D8A_7D5B_7D2E_7D00_7CCE_7C93;
    defparam RAM_inst1.INIT_A = 256'h82D4_8266_81FC_819E_8154_8123_810C_810F_8128_8150_817E_81AA_81CA_81D7_81CB_81A4;
    defparam RAM_inst1.INIT_B = 256'h8403_83F6_83E6_83DA_83D6_83DC_83EB_8402_841B_842F_8439_8432_8416_83E3_8399_833D;
    defparam RAM_inst1.INIT_C = 256'h7E9C_7EE5_7F30_7F83_7FE5_8055_80D3_815A_81E5_826B_82E6_834F_83A1_83DA_83FB_8407;
    defparam RAM_inst1.INIT_D = 256'h744C_7499_7500_7585_762B_76EF_77CC_78BA_79AD_7A9B_7B7A_7C42_7CEE_7D7C_7DEF_7E4D;
    defparam RAM_inst1.INIT_E = 256'h70D9_7044_6FE3_6FBB_6FCA_700A_7072_70F4_7182_720F_7290_72FF_7359_739F_73D9_7410;
    defparam RAM_inst1.INIT_F = 256'h753B_74FC_74F0_750E_7549_7590_75D1_75FA_75FE_75D1_7570_74DE_7424_734E_726E_7196;

endmodule

